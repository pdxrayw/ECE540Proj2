//	bot_if.v - Register interface to the Rojobot external world picoblaze 
//  Crystal Roberts
//  Ray Williams
//	
//	8-bit registers:
//			Loc_X		O	X (column) coordinate of Rojobot's current location
//			Loc_y		O 	Y (row) coordinate of Rojobot's current location
//			Sensors		O	Sensor values.  Rojobot contains a proximity sensor (left and right)
//						 	A proximity sensor is set to 1 if Rojobot detects an object in
//						  	front of it.  It also contains a black line sensor (left, center
//						  	and right).  Each black line sensor is set to 0 if there is
//							a black line under it and set to 1 if there is not black line
//							under it.
//			BotInfo		O 	Information on rojobot's current orientation and movement
//
//////////

module nexys4_bot_if(
	// interface to the picoblaze
	input 				Wr_Strobe,		// Write strobe - asserted to write I/O data
		 				Rd_Strobe,		// Read strobe - asserted to read I/O data
	input 		[7:0] 	AddrIn,			// I/O port address port_id
	input 		[7:0] 	DataIn,			// Data to be written to I/O register out_port
	output reg	[7:0] 	DataOut,		// I/O register data to picoblaze in_port

	// interface to the system	
	output reg 	[7:0]	MotCtl,			// (Port 0) Motor control input	into botsim
	input    	[7:0] 	LocX,			// (Port 1) X-coordinate of rojobot's location		
						LocY,			// (Port 2) Y-coordinate of rojobot's location
						BotInfo,		// (Port 3) Rojobot orientation and movement
						Sensors,		// (Port 4) Sensor readings
												
	// interface to the world map logic
//	output reg	[7:0]	MapX,			// (Port 8) Column address of world map location
//	output reg	[7:0]	MapY,			// (Port 9) Row address of world map location
//	input 		[1:0]	MapVal,			// (Port 10) Map value for location [row_addr, col_addr]	

	input               interrupt_ack,
	input				clk,			// system clock
						reset,			// system reset
	input   			upd_sysregs,	// flag from PicoBlaze to indicate that the system registers 
										// (LocX, LocY, Sensors, BotInfo)have been updated	
    input       [5:0]   db_btns,
    input       [15:0]  db_sw,
    output reg [15:0]   led, //out led
    output reg [4:0]    dig7, dig6, dig5, dig4, dig3, dig2, dig1, dig0, //7 seg display to sevenseg.v
    output reg [7:0]    dp,  //decimal point out to sevenseg.v   
    output reg          interrupt
		
);

// internal variables		
// used sot synchronize the register transfer so Application gets a consistant snapshot of the BOT status	
reg			load_sys_regs,			// Load system register flip-flop			
			load_dist_regs;			// Load distance register flip-flop
//reg         up_sys_reg = 0;

// holding registers for bot.  We want all registers to be updated
// at the same time (from system's point of view) to make sure
// the bot movement is consistent.
reg	[7:0] 	DataOut_int,					
            MotCtl_int,
            dp_int;
reg [15:0]   led_int;
reg [4:0]    dig7_int, dig6_int, dig5_int, dig4_int, dig3_int, dig2_int, dig1_int, dig0_int;
//reg          interrupt_int;
// read registers
always @(posedge clk) 
begin
    case(AddrIn[7:0])
    8'b0000_0000 : //pushbuttons inputs
    begin
    // format is: output(for this file) <= input (for this file)
    //dbbtns is total of [5:0]
        //dataout is to picoblaze
        DataOut[4:0] <= db_btns[5:1];
    end
    8'b0000_0001 : //slide switches
    begin
        DataOut <= db_sw[7:0];
    end
    8'b0000_1010 :// X coordinate of rojobot location
    begin
        DataOut <= LocX;
    end
    8'b0000_1011 : //(i))Y coordinate of rojobot location
    begin
        DataOut <= LocY;
    end
    8'b0000_1100 : //(i) Rojobot info register
    begin
        DataOut <= BotInfo;
    end
    8'b0000_1101 : //(i) Sensor register
    begin
        DataOut <= Sensors;
    end
    8'b0001_0000 : //(i) pushbutton inputs alternate port address
    begin
        DataOut[4:0] <= db_btns[5:1];
    end
    8'b0001_0001 : //(i) slide switches 15:8 (high byte of switches
    begin
        DataOut <= db_sw[15:8];
    end
    8'b0001_1010 : //(i) X coordinate of rojobot location
    begin
        DataOut <= LocX;
    end
    8'b0001_1011 : //(i) Y coordinate of rojobot location
    begin
        DataOut <= LocY;
    end
    8'b0001_1100 : //(i) Rojobot info register
    begin
        DataOut <= BotInfo;
    end
    8'b0001_1101 : //(i) Sensor register
    begin
        DataOut <= Sensors;
    end
    default : 
    begin
        DataOut <= 8'bXXXXXXXX;
    end
    endcase
end //always read registers


// write registers
always @(posedge clk) begin
	if (reset) begin

	end
	else begin
    if(Wr_Strobe) begin
    case (AddrIn[7:0])
    8'b0000_0010 : //(o) LEDs
        begin
        // format is: output(for this file) <= input (for this file)
        led[7:0] <= DataIn; //Datain is from picoblaze
        end
    8'b0000_0011 : // (o) digit 3 port address
        begin
        dig3 <= DataIn;
        end
    8'b0000_0100 : //(o) digit 2 port address
        begin
        dig2 <= DataIn;
        end
    8'b0000_0101 : //(o) digit 1 port address
        begin
        dig1 <= DataIn;
        end
    8'b0000_0110 : //(o) digit 0 port address
        begin
        dig0 <= DataIn;
        end
    8'b0000_0111 : //(o) decimal points 3:0 port address
        begin
        dp[3:0] <= DataIn[3:0];
        end
    8'b0000_1001 : //(o) Rojobot motor control output from system
        begin
        MotCtl <= DataIn;
        end
    8'b0001_0010 : //(o) LEDs 15:8 (high byte of switches)
        begin
        led[15:8] <= DataIn;
        end
    8'b0001_0011 : //(o) digit 7 port address
        begin
        dig7 <= DataIn;
        end
    8'b0001_0100 : //(o) digit 6 port address
        begin
        dig6 <= DataIn;
        end
    8'b0001_0101 : //(o) digit 5 port address
        begin
        dig5 <= DataIn;
        end
    8'b0001_0110 : //(o) digit 4 port address
        begin
        dig4 <= DataIn;
        end 
    8'b0001_0111 : //(o) decimal points 7:4 port address
        begin
        dp[7:4] <= DataIn; 
        end         
    8'b0001_1001 : //(o) Rojobot motor control output from system
        begin
        MotCtl <= DataIn; 
        end
    default :
        begin
        ;
        end
    endcase
    end
	end
end // always - write registers

	
always @ (posedge clk)
  begin
      if (interrupt_ack == 1'b1) begin
         interrupt <= 1'b0;
      end
      else if (upd_sysregs == 1'b1) begin
          interrupt <= 1'b1;
      end
      else begin
          interrupt <= interrupt;
      end
  end

endmodule
		
				

